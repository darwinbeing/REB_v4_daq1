-------------------------------------------------------------------------------
-- Title         : Version File
-- Project       : 
-------------------------------------------------------------------------------
-- File          : 
-- Author        : 
-- Created       : 
-------------------------------------------------------------------------------
-- Description:
-- Version Constant Module.
-------------------------------------------------------------------------------
-- Copyright (c) 2010 by SLAC National Accelerator Laboratory. All rights reserved.
-------------------------------------------------------------------------------
-- Modification history:
-- 
-------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

package Version is
-------------------------------------------------------------------------------
-- Version History
-------------------------------------------------------------------------------
  -- 00000001 Porting REB_v3 project under SLAC build system

  constant FPGA_VERSION_C : std_logic_vector(31 downto 0) := x"102c4005"; -- MAKE_VERSION

constant BUILD_STAMP_C : string := "REB_v4_top: Vivado v2015.3 (x86_64) Built Wed Oct 19 12:31:58 PDT 2016 by srusso";

end Version;

-------------------------------------------------------------------------------
-- Revision History:
-- 
-------------------------------------------------------------------------------
